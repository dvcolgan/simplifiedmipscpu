library ieee;
use ieee.std_logic_1164.all;

use work.mux4to1;

entity mux4to1_tb is
end mux4to1_tb;

architecture behavior of mux4to1_tb is
	component mux4to1
		port (S: in std_logic_vector(1 downto 0);
		      R: in std_logic_vector(3 downto 0);
		      O: out std_logic);
	end component;

	signal S: std_logic_vector(1 downto 0);
	signal R: std_logic_vector(3 downto 0);
	signal O: std_logic;
begin
	mux4to1_0: mux4to1 port map (S, R, O);

	process
		type pattern_type is record
			S0, S1, R0, R1, R2, R3: std_logic;
			O: std_logic;
		end record;

	type pattern_array is array (natural range <>) of pattern_type;
	constant patterns : pattern_array :=
		-- S0  S1   R0  R1  R2  R3   O
		(('0','0', '0','0','0','0', '0'),
		 ('0','0', '0','0','0','1', '0'),
		 ('0','0', '0','0','1','0', '0'),
		 ('0','0', '0','0','1','1', '0'),
		 ('0','0', '0','1','0','0', '0'),
		 ('0','0', '0','1','0','1', '0'),
		 ('0','0', '0','1','1','0', '0'),
		 ('0','0', '0','1','1','1', '0'),
		 ('0','0', '1','0','0','0', '1'),
		 ('0','0', '1','0','0','1', '1'),
		 ('0','0', '1','0','1','0', '1'),
		 ('0','0', '1','0','1','1', '1'),
		 ('0','0', '1','1','0','0', '1'),
		 ('0','0', '1','1','0','1', '1'),
		 ('0','0', '1','1','1','0', '1'),
		 ('0','0', '1','1','1','1', '1'),

		 ('0','1', '0','0','0','0', '0'),
		 ('0','1', '0','0','0','1', '0'),
		 ('0','1', '0','0','1','0', '1'),
		 ('0','1', '0','0','1','1', '1'),
		 ('0','1', '0','1','0','0', '0'),
		 ('0','1', '0','1','0','1', '0'),
		 ('0','1', '0','1','1','0', '1'),
		 ('0','1', '0','1','1','1', '1'),
		 ('0','1', '1','0','0','0', '0'),
		 ('0','1', '1','0','0','1', '0'),
		 ('0','1', '1','0','1','0', '1'),
		 ('0','1', '1','0','1','1', '1'),
		 ('0','1', '1','1','0','0', '0'),
		 ('0','1', '1','1','0','1', '0'),
		 ('0','1', '1','1','1','0', '1'),
		 ('0','1', '1','1','1','1', '1'),

		 ('1','0', '0','0','0','0', '0'),
		 ('1','0', '0','0','0','1', '0'),
		 ('1','0', '0','0','1','0', '0'),
		 ('1','0', '0','0','1','1', '0'),
		 ('1','0', '0','1','0','0', '1'),
		 ('1','0', '0','1','0','1', '1'),
		 ('1','0', '0','1','1','0', '1'),
		 ('1','0', '0','1','1','1', '1'),
		 ('1','0', '1','0','0','0', '0'),
		 ('1','0', '1','0','0','1', '0'),
		 ('1','0', '1','0','1','0', '0'),
		 ('1','0', '1','0','1','1', '0'),
		 ('1','0', '1','1','0','0', '1'),
		 ('1','0', '1','1','0','1', '1'),
		 ('1','0', '1','1','1','0', '1'),
		 ('1','0', '1','1','1','1', '1'),

		 ('1','1', '0','0','0','0', '0'),
		 ('1','1', '0','0','0','1', '1'),
		 ('1','1', '0','0','1','0', '0'),
		 ('1','1', '0','0','1','1', '1'),
		 ('1','1', '0','1','0','0', '0'),
		 ('1','1', '0','1','0','1', '1'),
		 ('1','1', '0','1','1','0', '0'),
		 ('1','1', '0','1','1','1', '1'),
		 ('1','1', '1','0','0','0', '0'),
		 ('1','1', '1','0','0','1', '1'),
		 ('1','1', '1','0','1','0', '0'),
		 ('1','1', '1','0','1','1', '1'),
		 ('1','1', '1','1','0','0', '0'),
		 ('1','1', '1','1','0','1', '1'),
		 ('1','1', '1','1','1','0', '0'),
		 ('1','1', '1','1','1','1', '1'));

	begin
		assert false report "Testing mux4to1" severity note;
		for c in patterns'range loop
			S(0) <= patterns(c).S0;
			S(1) <= patterns(c).S1;
			R(0) <= patterns(c).R0;
			R(1) <= patterns(c).R1;
			R(2) <= patterns(c).R2;
			R(3) <= patterns(c).R3;
			wait for 1 ns;
			assert O = patterns(c).O
				report "test failed" severity error;
		end loop;

		wait;
	end process;
end behavior;

