library ieee;
use ieee.std_logic_1164.all;

use work.mux32x32to1;
use work.datatypes.bus32x32;

entity mux32x32to1_tb is
end mux32x32to1_tb;

architecture behavior of mux32x32to1_tb is
	component mux32x32to1
		port (S: in std_logic_vector(4 downto 0);
		      R: in bus32x32;
		      O: out std_logic_vector(31 downto 0));
	end component;

	signal S: std_logic_vector(4 downto 0);
	signal R: bus32x32;
	signal O: std_logic_vector(31 downto 0);
begin
	mux32x32to1_0: mux32x32to1 port map (S, R, O);

	process
	begin
		assert false report "Testing mux32x32to1" severity note;
		R(0) <= X"0000_0000";
		R(1) <= X"0000_1111";
		R(2) <= X"0000_2222";
		R(3) <= X"0000_3333";
		R(4) <= X"0000_4444";
		R(5) <= X"0000_5555";
		R(6) <= X"0000_6666";
		R(7) <= X"0000_7777";
		R(8) <= X"0000_8888";
		R(9) <= X"0000_9999";
		R(10) <= X"0000_AAAA";
		R(11) <= X"0000_BBBB";
		R(12) <= X"0000_CCCC";
		R(13) <= X"0000_DDDD";
		R(14) <= X"0000_EEEE";
		R(15) <= X"0000_FFFF";
		R(16) <= X"1111_0000";
		R(17) <= X"2222_0000";
		R(18) <= X"3333_0000";
		R(19) <= X"4444_0000";
		R(20) <= X"5555_0000";
		R(21) <= X"6666_0000";
		R(22) <= X"7777_0000";
		R(23) <= X"8888_0000";
		R(24) <= X"9999_0000";
		R(25) <= X"AAAA_0000";
		R(26) <= X"BBBB_0000";
		R(27) <= X"CCCC_0000";
		R(28) <= X"DDDD_0000";
		R(29) <= X"EEEE_0000";
		R(30) <= X"FFFF_0000";
		R(31) <= X"FFFF_FFFF";
		S <= "00000";
		wait for 1 ns;
		assert O = X"0000_0000" report "test failed" severity error;
		S <= "00001";
		wait for 1 ns;
		assert O = X"0000_1111" report "test failed" severity error;
		S <= "00010";
		wait for 1 ns;
		assert O = X"0000_2222" report "test failed" severity error;
		S <= "00011";
		wait for 1 ns;
		assert O = X"0000_3333" report "test failed" severity error;
		S <= "00100";
		wait for 1 ns;
		assert O = X"0000_4444" report "test failed" severity error;
		S <= "00101";
		wait for 1 ns;
		assert O = X"0000_5555" report "test failed" severity error;
		S <= "00110";
		wait for 1 ns;
		assert O = X"0000_6666" report "test failed" severity error;
		S <= "00111";
		wait for 1 ns;
		assert O = X"0000_7777" report "test failed" severity error;
		S <= "01000";
		wait for 1 ns;
		assert O = X"0000_8888" report "test failed" severity error;
		S <= "01001";
		wait for 1 ns;
		assert O = X"0000_9999" report "test failed" severity error;
		S <= "01010";
		wait for 1 ns;
		assert O = X"0000_AAAA" report "test failed" severity error;
		S <= "01011";
		wait for 1 ns;
		assert O = X"0000_BBBB" report "test failed" severity error;
		S <= "01100";
		wait for 1 ns;
		assert O = X"0000_CCCC" report "test failed" severity error;
		S <= "01101";
		wait for 1 ns;
		assert O = X"0000_DDDD" report "test failed" severity error;
		S <= "01110";
		wait for 1 ns;
		assert O = X"0000_EEEE" report "test failed" severity error;
		S <= "01111";
		wait for 1 ns;
		assert O = X"0000_FFFF" report "test failed" severity error;
		S <= "10000";
		wait for 1 ns;
		assert O = X"1111_0000" report "test failed" severity error;
		S <= "10001";
		wait for 1 ns;
		assert O = X"2222_0000" report "test failed" severity error;
		S <= "10010";
		wait for 1 ns;
		assert O = X"3333_0000" report "test failed" severity error;
		S <= "10011";
		wait for 1 ns;
		assert O = X"4444_0000" report "test failed" severity error;
		S <= "10100";
		wait for 1 ns;
		assert O = X"5555_0000" report "test failed" severity error;
		S <= "10101";
		wait for 1 ns;
		assert O = X"6666_0000" report "test failed" severity error;
		S <= "10110";
		wait for 1 ns;
		assert O = X"7777_0000" report "test failed" severity error;
		S <= "10111";
		wait for 1 ns;
		assert O = X"8888_0000" report "test failed" severity error;
		S <= "11000";
		wait for 1 ns;
		assert O = X"9999_0000" report "test failed" severity error;
		S <= "11001";
		wait for 1 ns;
		assert O = X"AAAA_0000" report "test failed" severity error;
		S <= "11010";
		wait for 1 ns;
		assert O = X"BBBB_0000" report "test failed" severity error;
		S <= "11011";
		wait for 1 ns;
		assert O = X"CCCC_0000" report "test failed" severity error;
		S <= "11100";
		wait for 1 ns;
		assert O = X"DDDD_0000" report "test failed" severity error;
		S <= "11101";
		wait for 1 ns;
		assert O = X"EEEE_0000" report "test failed" severity error;
		S <= "11110";
		wait for 1 ns;
		assert O = X"FFFF_0000" report "test failed" severity error;
		S <= "11111";
		wait for 1 ns;
		assert O = X"FFFF_FFFF" report "test failed" severity error;

		wait;
	end process;
end behavior;

